`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Lafayette College
// Engineer: John Nestor
//
// Create Date: 01/10/2019 10:03:33 AM
// Design Name: BRAM storage for adafruit LED matrix
// Module Name: pixel_ram
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module pixel_ram(
  input logic        clk,
  input logic        rst,
  input logic [12:0] rdaddr_pix_upper,
  output logic [3:0] dout_pix_upper,
  input logic [12:0] rdaddr_pix_lower,
  output logic [3:0] dout_pix_lower,
  input logic        we_lower,
  input logic [9:0]  wraddr_col_lower,
  input logic [31:0] din_col_lower
  );

  logic [3:0] we_lower_byte;  // byte write enable
  assign we_lower_byte = { 4 {we_lower} };

  // Upper RAM (read-only)
  BRAM_SDP_MACRO #(
  .BRAM_SIZE("36Kb"), // Target BRAM, "18Kb" or "36Kb"
  .DEVICE("7SERIES"), // Target device: "7SERIES"
  .WRITE_WIDTH(32),    // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
  .READ_WIDTH(4),     // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
  .DO_REG(0),         // Optional output register (0 or 1)
  .INIT_FILE ("NONE"),
  .SIM_COLLISION_CHECK ("ALL"), // Collision check enable "ALL", "WARNING_ONLY",
  //   "GENERATE_X_ONLY" or "NONE"
  .SRVAL(72'h000000000000000000), // Set/Reset value for port output
  .INIT(72'h000000000000000000),  // Initial values on output port
  .WRITE_MODE("WRITE_FIRST"),  // Specify "READ_FIRST" for same clock or synchronous clocks
  //   Specify "WRITE_FIRST for asynchronous clocks on ports

  .INIT_00(256'h11111111_00000000_00000000_44444444_00000004_00000004_00000004_22222222),
.INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_20 (256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_21212121),
.INIT_21 (256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
.INIT_22 (256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
.INIT_23 (256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
.INIT_24 (256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
.INIT_25 (256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
.INIT_26 (256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
.INIT_27 (256'h20000021_20000021_20000021_21212121_00000000_00000000_00000000_00000000),
.INIT_28 (256'h00000000_00000020_00000001_00000001_00000001_21212120_00000000_20000021),
.INIT_29 (256'h00000000_00000000_00000000_20000021_20000021_20000021_20000021_21212121),
.INIT_2A (256'h00010000_00010000_00010000_00010000_00000000_00000000_00000000_00000000),
.INIT_2B (256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00010000),
.INIT_2C (256'h00000000_00000000_00000000_00000001_20000001_01000001_00200001_00012120),
.INIT_2D (256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
.INIT_2E (256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
.INIT_2F (256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
.INIT_30 (256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
.INIT_31 (256'h00000000_21212120_20000001_20000001_20000001_00000001_00000000_00000000),
.INIT_32 (256'h20000001_00000001_00000000_21212121_00000021_00000021_00000021_21212121),
.INIT_33 (256'h20000001_20000001_00000001_00000120_00000000_21212120_20000001_20000001),
.INIT_34 (256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_01212120)
  /*
  .INIT_04(256'h10000004_01226640_00000000_10000004_10006004_10006004_10006004_11226644),
  .INIT_05(256'h10006004_10006004_10006004_11226644_00000000_01000040_10000004_10000004),
  .INIT_06(256'h10020004_10200004_11000040_00000000_00000000_00000000_00000000_10000004),
  .INIT_07(256'h11000040_00000000_10000000_11226644_10000040_00000000_10000640_10006004),
  .INIT_08(256'h00000000_00000000_00000000_00000000_10000640_10006004_10020004_10200004)*/
  // everything else is blank!

  ) BRAM_UPPER (
  .DO(dout_pix_upper),         // Output read data port, width defined by READ_WIDTH parameter
  .DI(32'd0),         // Input write data port, width defined by WRITE_WIDTH parameter
  .RDADDR(rdaddr_pix_upper), // Input read address, width defined by read port depth
  .RDCLK(clk),   // 1-bit input read clock
  .RDEN(1'b1),     // 1-bit input read port enable
  .REGCE(1'b0),   // 1-bit input read output register enable
  .RST(rst),       // 1-bit input reset
  .WE(4'b0000),         // Input write enable, width defined by write port depth
  .WRADDR(10'd0), // Input write address, width defined by write port depth
  .WRCLK(clk),   // 1-bit input write clock
  .WREN(1'b1)      // 1-bit input write port enable
  );

  // Lower half-matrix RAM
  BRAM_SDP_MACRO #(
  .BRAM_SIZE("36Kb"), // Target BRAM, "18Kb" or "36Kb"
  .DEVICE("7SERIES"), // Target device: "7SERIES"
  .WRITE_WIDTH(32),    // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
  .READ_WIDTH(4),     // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
  .DO_REG(0),         // Optional output register (0 or 1)
  .INIT_FILE ("NONE"),
  .SIM_COLLISION_CHECK ("ALL"), // Collision check enable "ALL", "WARNING_ONLY",
  //   "GENERATE_X_ONLY" or "NONE"
  .SRVAL(72'h000000000000000000), // Set/Reset value for port output
  .INIT(72'h000000000000000000),  // Initial values on output port
  .WRITE_MODE("WRITE_FIRST"),  // Specify "READ_FIRST" for same clock or synchronous clocks
  //   Specify "WRITE_FIRST for asynchronous clocks on ports
  .INIT_00(256'h11111111_00000000_00000000_44444444_40000000_00000004_40000000_22222222),
.INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_10 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_11 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_12 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_13 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_14 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_15 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_16 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_17 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_18 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_19 (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1A (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1B (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1C (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1D (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1E (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_1F (256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_20 (256'h20010100_01200000_00000000_20000000_20000000_20000000_20000000_21212121),
.INIT_21 (256'h00000020_00010020_21212100_00010000_00000000_01202000_20010100_20010100),
.INIT_22 (256'h00000000_01202000_20010100_20010100_20010100_01200000_00000000_00000100),
.INIT_23 (256'h20202000_01210000_00000000_01212000_20200000_20200000_20200000_00012000),
.INIT_24 (256'h20002000_21212120_00002000_00000000_00000000_00210000_20202000_20202000),
.INIT_25 (256'h00000000_01000000_20002000_21212120_00002000_00000000_00000000_01000000),
.INIT_26 (256'h00000000_00000000_00000000_00210000_20202000_20202000_20202000_01210000),
.INIT_27 (256'h21000001_21000001_21000001_21212121_00000000_00000000_00000000_00000000),
.INIT_28 (256'h00000000_01000000_20000000_20000000_20000000_01212121_00000000_21000001),
.INIT_29 (256'h00000000_00000000_00000000_21000001_21000001_21000001_21000001_21212121),
.INIT_2A (256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
.INIT_2B (256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
.INIT_2C (256'h20000000_01212000_00000000_01212121_20000000_20000000_20000000_20000000),
.INIT_2D (256'h00002000_21210000_00002000_21212000_00000000_21212000_01000000_20000000),
.INIT_2E (256'h00000000_21210000_00002000_21210000_00002000_21212000_00000000_21210000),
.INIT_2F (256'h00010000_21212000_00000000_00210000_20202000_20202000_20202000_01210000),
.INIT_30 (256'h00000000_00000000_00000000_00000000_00000000_00210000_00002000_00002000),
.INIT_31 (256'h00000000_20000000_20000000_20000000_20000000_01212121_00000000_00000000),
.INIT_32 (256'h20000000_01212121_00000000_21212121_21000000_21000000_21000000_21212121),
.INIT_33 (256'h20000000_20000000_20000000_01200000_00000000_20000000_20000000_20000000),
.INIT_34 (256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_01212121)
  // everything else is blank!

  ) BRAM_LOWER (
  .DO(dout_pix_lower),         // Output read data port, width defined by READ_WIDTH parameter
  .DI(din_col_lower),         // Input write data port, width defined by WRITE_WIDTH parameter
  .RDADDR(rdaddr_pix_lower), // Input read address, width defined by read port depth
  .RDCLK(clk),   // 1-bit input read clock
  .RDEN(1'b1),     // 1-bit input read port enable
  .REGCE(1'b0),   // 1-bit input read output register enable
  .RST(rst),       // 1-bit input reset
  .WE(we_lower_byte),         // Input write enable, width defined by write port depth
  .WRADDR(wraddr_col_lower), // Input write address, width defined by write port depth
  .WRCLK(clk),   // 1-bit input write clock
  .WREN(1'b1)      // 1-bit input write port enable
  );

endmodule
